library verilog;
use verilog.vl_types.all;
entity DividerTest is
end DividerTest;

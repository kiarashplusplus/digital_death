library verilog;
use verilog.vl_types.all;
entity gcd_test is
end gcd_test;

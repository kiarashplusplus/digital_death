library verilog;
use verilog.vl_types.all;
entity SirenTest is
end SirenTest;
